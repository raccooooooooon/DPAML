DIM
FREQ GHZ
LNG MM
CAP PF
IND NH
RES OH

CKT
MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
MLIN 1 0 W=1.52 L=33.42
DEF1P 1 SHORT2
RES 2 3 R=1.42
IND 3 4 L=5.1
CAP 4 0 C=0.83
DEF1P 2 CIR1

OUT
SHORT2 MAG[Y1] GR1
SHORT2 IM[Y1] GR2
SHORT2 S11
CIR1 MAG[Y1] GR1
CIR1 IM[Y1] GR2

FREQ
SWEEP 2 3 0.005

GRID
GR1 0 0.8 0.1
GR2 -0.5 0.5 0.1
 
 