! Basic CKT file

DIM
   FREQ  MHZ
   RES  OH
   LNG  MM
   ANG DEG
   IND NH
   CAP PF

CKT
   MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=1.52 L=5
   MLIN 2 3 W=1.52 L=9.83
   MLIN 2 4 W=1.52 L=2.94
   MLOC 3 W=1.52 L=0
   RES 4 0 R=15
   !IND 5 0 L=0.8
   DEF1P 1 EXP2

OUT
   EXP2 DB[S11] GR1

FREQ
   SWEEP 1000 4000 10

GRID
   RANGE 1000 4000 100
   GR1 -40 0 5
 
 
 
 