/*******************************************************************************************************************
* �ɮצW�١Ghw01_7seg.v
* �ҲզW�١G�C�q��ܸѽX��
* �\    ��G�N4bits�G�i��Ʀr�ର�@�C�q��ܾ��A�åH�Q���i����ܡC
* ��J�ѼơGdin		4bits�G�i��Ʀr           
* ��X�ѼơGdout	7bits�C�q��ܾ���J�}
* ��    ���G�C�q��ܾ����@�����A�G�T��0���G�C
													JH design
*******************************************************************************************************************/


module hw01_7seg(din,dout); 
input 	[3:0]	din;
output	[6:0]	dout;
reg		[6:0]	dout;
always@(din)
begin
	case(din)
	 	4'b0000:dout<=7'b1000000;
	 	4'b0001:dout<=7'b1111001;
	 	4'b0010:dout<=7'b0100100;
	 	4'b0011:dout<=7'b0110000;
	 	4'b0100:dout<=7'b0011001;
	 	4'b0101:dout<=7'b0010010;
	 	4'b0110:dout<=7'b0000010;
	 	4'b0111:dout<=7'b1111000;
		4'b1000:dout<=7'b0000000;
	 	/*�Цb�����g�{���X�A�ϵ{���X����*/
	endcase
end
endmodule
