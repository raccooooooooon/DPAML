DIM
FREQ MHZ
RES OH
LNG MM
ANG DEG
IND NH
CAP PF

CKT
MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
IND 1 2 L=10.212
CAP 2 0 C=0.803
RES 2 3 R=240
IND 3 0 L=12
DEF1P 1 EXP1

MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
CAP 1 2 C=0.766
IND 2 0 L=16.056
RES 2 3 R=240
IND 3 0 L=12
DEF1P 1 EXP2

FREQ
SWEEP 0 3000 10

OUT
EXP1 DB[S11] GR1
EXP2 DB[S11] GR2

GRID
GR1 -60 0 5
GR2 -60 0 5
 