DIM
FREQ GHZ
LNG MM
CAP PF
IND NH
RES OH

CKT
MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
MLIN 1 0 W=1.52 L=16.71
DEF1P 1 short4
RES 2 0 R=3520.26
IND 2 0 L=4.14
CAP 2 0 C=1.02
DEF1P 2 CIR1

OUT
short4 MAG[Z1] GR1
short4 IM[Z1] GR2
short4 S11
CIR1 MAG[Z1] GR1
CIR1 IM[Z1] GR2

FREQ
SWEEP 2 3 0.005

GRID
GR1 0 4000 500
GR2 -2000 2000 500
 
 
 
 