DIM
FREQ GHZ
LNG MM
CAP PF
IND NH
RES OH

CKT
MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
MLIN 1 2 W=1.52 L=16.71
DEF1P 1 open4
RES 3 4 R=0.71
IND 4 5 L=2.55
CAP 5 0 C=1.65
DEF1P 3 CIR1

OUT
open4 MAG[Y1] GR1
open4 IM[Y1] GR2
open4 S11
CIR1 MAG[Y1] GR1
CIR1 IM[Y1] GR2

FREQ
SWEEP 2 3 0.005

GRID
GR1 0 1.5 0.3
GR2 -1 1 0.2
 
 
 
 
 
 