


module tb;



endmodule
