DIM
  LNG M
  FREQ GHZ
  IND NH
  CAP PF
  RES OH
  ANG DEG

VAR
  L1=1197.3
  C1=9.28
  ZTL=359.193
  ETL=120
  FRE=1
  LINE=0.1

EQN
  LAT=L1*LINE/4
  CAT=C1*LINE/2
  LATK=L1*LINE/2000
  CATK=C1*LINE/1000
  LAP=L1*LINE/2
  CAP=C1*LINE/4
  LAPK=L1*LINE/1000
  CAPK=C1*LINE/2000

CKT 
  TLIN 1 2 Z^ZTL E^ETL F^FRE
  RES 2 0 R=50
  DEF1P 1  EXP1
!
  IND 3 4 L^LAT
  IND 4 5 L^LAT
  CAP 4 0 C^CAT
  DEF2P 3 5 LCCELL
  LCCELL 6  7
  LCCELL 7  8
  RES 8 0 R=50
  DEF1P 6 LC1
!
  IND 9 10  L^LATK
  IND 10 11 L^LATK
  CAP 10 0  C^CATK
  DEF2P 9 11 CELL1
  CELL1 12 13
  CELL1 13 14
  CELL1 14 15
  CELL1 15 16
  CELL1 16 17
  DEF2P 12 17 CELL5
  CELL5 18 19
  CELL5 19 20
  CELL5 20 21
  CELL5 21 22
  CELL5 22 23
  DEF2P 18 23 CELL25
  CELL25 24 25
  CELL25 25 26
  CELL25 26 27
  CELL25 27 28
  CELL25 28 29
  CELL25 29 30
  CELL25 30 31
  CELL25 31 32
  DEF2P 24 32 CELL200
  CELL200 33 34
  CELL200 34 35
  CELL200 35 36
  CELL200 36 37
  CELL200 37 38
  RES 38 0 R=50
  DEF1P 33 LC2
!
OUT
  EXP1 DB[S11] GR1
  EXP1 RE[Z1] GR2
  EXP1 IM[Z1] GR3
  LC1 DB[S11] GR1
  LC1 RE[Z1] GR2
  LC1 IM[Z1] GR3
  LC2 DB[S11] GR1
  LC2 RE[Z1] GR2
  LC2 IM[Z1] GR3

FREQ
  SWEEP 0 2 0.005

GRID
  GR1 -50 5 5
  GR2 0 3000 500
  GR3 -2000 2000 500
 
 