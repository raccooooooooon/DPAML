DIM
   FREQ  MHZ
   RES  OH
   LNG  MM
   ANG DEG
   IND NH
   CAP PF

CKT
   MSUB ER=4.7 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=5.33541 L=70
   DEF1P 1 EXP1

FREQ
   SWEEP 1000 4000 50
OUT
   EXP1  DB[S11] GR1 
   EXP1  MAG[z1] GR2
GRID
   RANGE 1000 4000 50
   GR1 -5 0 5
   GR2 0 300 10