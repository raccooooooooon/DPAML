DIM
FREQ GHZ
LNG MM
CAP PF
IND NH
RES OH

CKT
MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.02
MLIN 1 2 W=1.52 L=33.42
DEF1P 1 open2
RES 3 0 R=1760.13
IND 3 0 L=2.07
CAP 3 0 C=2.04
DEF1P 3 CIR1

OUT
open2 MAG[Z1] GR1
open2 IM[Z1] GR2
open2 S11
CIR1 MAG[Z1] GR1
CIR1 IM[Z1] GR2

FREQ
SWEEP 2 3 0.005

GRID
GR1 0 2000 500
GR2 -1000 1000 500
 
 
 
 
 