DIM
   FREQ  GHZ
   RES   OH
   LNG   MM
   ANG   DEG
   IND   NH
   CAP   PF

CKT
   MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 0 W=1.52 L=6
   MLIN 1 2 W=1.52 L=0.85
   RES 2 3 R=22.5
   CAP 3 0 C=1.768
   DEF1P 1 CIR1

OUT
   CIR1 DB[S11] GR1

FREQ
   SWEEP 2 4 0.005

GRID
   GR1 0 -60 5
 
 
 
 
 