DIM
  LNG M
  FREQ GHZ
  IND NH
  CAP PF
  RES OH
  ANG DEG

VAR
  L1=1197.3
  C1=4.64
  ZTL=359.193
  ETL=120
  FRE=1
  LINE=0.1

EQN
  LA=L1*LINE/2
  CA=C1*LINE/2
  LA1=L1*LINE/1000
  CA1=C1*LINE/1000
CKT 
  TLIN 1 2 Z^ZTL E^ETL F^FRE
  RES 2 0 R=50
  DEF1P 1  EXP1

  CAP 3 0 C^CA
  IND 3 4 L^LA
  CAP 4 0 C^CA
  DEF2P 3 4 LCCELL
  LCCELL 34 35
  LCCELL 35 36
  RES 36 0 R=50
  DEF1P 34 LC1

  CAP 5 0 C^CA1
  IND 5 6 L^LA1
  CAP 6 0 C^CA1
  DEF2P 5 6 CELL1
  CELL1 7 8
  CELL1 8 9
  CELL1 9 10
  CELL1 10 11
 CELL1 11 12
  DEF2P 7 12 CELL5
  CELL5 13 14
  CELL5 14 15
  CELL5 15 16
  CELL5 16 17
  CELL5 17 18
  DEF2P 13 18 CELL25

  CELL25 19 20
  CELL25 20 21
  CELL25 21 22
  CELL25 22 23
  CELL25 23 24
  CELL25 24 25
  CELL25 25 26
  CELL25 26 27
  DEF2P 19 27 CELL200

  CELL200 28 29
  CELL200 29 30
  CELL200 30 31
  CELL200 31 32
  CELL200 32 33
  RES 33 0 R=50
  DEF1P 28 LC2
OUT
  EXP1 DB[S11] GR1
  EXP1 RE[Z1] GR2
  EXP1 IM[Z1] GR3
  LC1 DB[S11] GR1
  LC1 RE[Z1] GR2
  LC1 IM[Z1] GR3
  LC2 DB[S11] GR1
  LC2 RE[Z1] GR2
  LC2 IM[Z1] GR3


FREQ
  SWEEP 0 2 0.005


GRID
  GR1 -50 5 5
  GR2 0 20000 1000
  GR3 -10000 10000 1000