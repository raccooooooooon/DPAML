DIM
  LNG M
  FREQ GHZ
  IND NH
  CAP PF
  RES OH
  ANG DEG

VAR
  L1=598.65
  C1=9.28
  ZTL=359.193
  ETL=120
  FRE=1
  LINE=0.1

EQN
  LA=L1*LINE/2
  CA=C1*LINE/2
  LA1=L1*LINE/1000
  CA1=C1*LINE/1000
CKT 
  TLIN 1 2 Z^ZTL E^ETL F^FRE
  RES 2 0 R=50
  DEF1P 1  EXP1

  IND 3 4 L^LA
  CAP 4 0 C^CA
  IND 4 5 L^LA
  DEF2P 3 5 LCCELL
  LCCELL 36 37
  LCCELL 37 38
  RES 38 0 R=50
  DEF1P 36 LC1

  IND 6 7 L^LA1
  CAP 7 0 C^CA1
  IND 7 8 L^LA1
  DEF2P 6  8  CELL1
  CELL1 9  10
  CELL1 10 11
  CELL1 11 12
  CELL1 12 13
  CELL1 13 14
  DEF2P 9 14 CELL5

  CELL5 15 16
  CELL5 16 17
  CELL5 17 18
  CELL5 18 19
  CELL5 19 20
  DEF2P 15 20 CELL25

  CELL25 21 22
  CELL25 22 23
  CELL25 23 24
  CELL25 24 25
  CELL25 25 26
  CELL25 26 27
  CELL25 27 28
  CELL25 28 29
  DEF2P 21 29 CELL200

  CELL200 30 31
  CELL200 31 32
  CELL200 32 33
  CELL200 33 34
  CELL200 34 35
  RES 35 0 R=50
  DEF1P 30 LC2
OUT
  EXP1 DB[S11] GR1
  EXP1 RE[Z1] GR2
  EXP1 IM[Z1] GR3
  LC1 DB[S11] GR1
  LC1 RE[Z1] GR2
  LC1 IM[Z1] GR3
  LC2 DB[S11] GR1
  LC2 RE[Z1] GR2
  LC2 IM[Z1] GR3


FREQ
  SWEEP 0 2 0.005


GRID
  GR1 -50 5 5
  GR2 0 3000 500
  GR3 -2000 2000 500