DIM
   FREQ  GHZ
   RES   OH
   LNG   MM
   ANG   DEG
   IND   NH
   CAP   PF
CKT
   MSUB ER=4.4 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=1.52 L=50
   DEF2P 1 2 L0.8

   MSUB ER=4.4 H=1.6 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 3 4 W=3.05 L=50
   DEF2P 3 4 L1.6
   
FREQ
   SWEEP 0 9 0.1

OUT
   L0.8 DB[S21] GR1
   L1.6 DB[S21] GR1

GRID
   RANGE 0 9 1
   GR1 -2.5 0.5 0.5
