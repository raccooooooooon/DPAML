DIM
   FREQ GHZ
   LNG MM
   ANG DEG
   RES OH
   CAP PF
   IND NH

CKT
   MSUB ER=4.7 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=3.14015 L=44.1985
   RES 2 0 R=27
   DEF1P 1 EXP312
   
   MSUB ER=4.7 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=2.3549 L=52.4905
   RES 2 0 R=27
   DEF1P 1 EXP314
   

FREQ
   SWEEP 0.1 3 0.01

OUT
   EXP312 MAG[Z1] GR1
   EXP312 DB[S11] GR2
   EXP314 MAG[Z1] GR3
   EXP314 DB[S11] GR4
	 

GRID
   GR1 0 50 10
   GR2 0 -15 5
   GR3 0 50 10
   GR4 0 -45 5
 