DIM
   FREQ MHZ
   RES  OH
   LNG  MM
   ANG  DEG

CKT
TLIN 1 2 Z=100 E=54.735 F=1000
TLSC 1 0 Z=100 E=54.61 F=1000
RES 2 0 R=200
DEF1P 1 MATCH

TERM
Z0=100
MATCH 0 0 0 0

OUT
MATCH DB[S11] GR1

FREQ
SWEEP 50 3000 50

GRID
RANGE 50 3000 50
GR1 -30 0 5
 