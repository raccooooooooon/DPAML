DIM
FREQ GHZ
LNG MM
CAP PF
IND NH
RES OH

CKT
IND 1 2 L=0.265
IND 1 0 L=2.411
RES 2 3 R=22.5
CAP 3 0 C=1.768
DEF1P 1 CIR1

OUT
CIR1 DB[S11] GR1

FREQ
SWEEP 2 4 0.005

GRID
GR1 0 -60 5
 
 
 
 
 