DIM
FREQ GHZ
RES OH
LNG MM
ANG DEG
IND NH
CAP PF

CKT
MSUB ER=4.7 H=0.8 T=0.01 RHO=0 RGH=0
TAND TAND=0.01
MLIN 1 2 W=2.35389 L=39.0465
RES 2 0 R=27
DEF1P 1 EXP1

FREQ
SWEEP 0 3 0.1

OUT
EXP1 DB[S11] GR1
EXP1 MAG[Z1] GR2

GRID
GR1 -50 0 5
GR2  0  60 10
 
 
 
 