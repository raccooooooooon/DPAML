DIM
FREQ	GHZ
RES	OH
LNG	MM
ANG	DEG
IND	NH
CAP	PF

CKT
MSUB	ER=4.7	H=0.8	T=0.035	RHO=0	RGH=0
TAND		TAND=0.02
MLIN	1	2	W=2.04411	L=70
RES	2	0	R=0
DEF1P	1	EXP1

FREQ
SWEEP	0	4	0.01

OUT
EXP1	DB[S11]	GR1
EXP1	MAG[z1]	GR2

GRID
RANGE	0	4	0.01
GR1	-2	0.5	0.01
GR2	-100	1500	100
 