DIM
   FREQ  MHZ
   RES  OH
   LNG  MM
   ANG DEG
   IND NH
   CAP PF

CKT
   MSUB ER=4.7 H=0.8 T=0.01 RHO=0 RGH=0
   TAND TAND=0.02
   MLIN 1 2 W=1.44584 L=29.5
   MLIN 2 0 W=1.44584 L=19.5861
   MLIN 2 4 W=1.44584 L=58.5649
   RES 4 5 R=27
   CAP 5 0 C=10
   DEF1P 1 EXP1

FREQ
   SWEEP 100 3000 10

OUT
   EXP1 DB[S11] GR1
   EXP1 MAG[Z1] GR2

GRID
   RANGE 100 3000 100
   GR1 -40 0 5 
   GR2 0 350 30